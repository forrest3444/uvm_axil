`timescale 1ns/1ps
`include "uvm_macros.svh"

import uvm_pkg::*;
`include "axil_drv.sv"

module top_tb;

