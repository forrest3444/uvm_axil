`ifndef AXIL_ENV__SV
`define AXIL_ENV__SV

class axil_env extends uvm_env;
	:
