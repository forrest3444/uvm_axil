`ifndef AXIL_AGENT__SV
`define AXIL_AGENT__SV

class axil_agent extends uvm_agent;
	axil_driver         drv;
	axil_:
