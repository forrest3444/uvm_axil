`ifndef	AXIL_SEQ__SV
`define AXIL_SEQ__SV

class :wq

